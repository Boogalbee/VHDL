library ieee;
use ieee.std_logic_1164.all;

entity my_xor is
	port(a,b,c: IN std_logic; f: OUT std_logic);
end my_xor;
architecture behav of my_xor is
begin
	f <= a XOR b XOR c;
end;
